///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: IITB
//
// File: and_gate.v
// Targeted device: <Family::ProASIC3E> <Die::A3PE1500> <Package::208 PQFP>
// Author: Abhijeet
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

module control_signal (miso,miso_probe,ss1,ss2);

input miso;
output reg miso_probe;
input ss1;
input ss2;
//and (y,a,b);

always @*
miso_probe <= miso;

endmodule

