///////////////////////////////////////////////////////////////////////////////////////////////////
// Company: IITB
//
// File: and_gate.v
// Targeted device: <Family::ProASIC3E> <Die::A3PE1500> <Package::208 PQFP>
// Author: Abhijeet
//
/////////////////////////////////////////////////////////////////////////////////////////////////// 

module control_signal (miso,ss1,ss2);

input miso;

output reg ss1;
output reg ss2;
//and (y,a,b);

endmodule

